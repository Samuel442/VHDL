
-- IMPLEMENTA��O DE UM CIRCUITO L�GICO COMBINACIONAL A PARTIR DA TABELA DA VERDADE 1 DO ARQUIVO ANEXO (COMPLEMENTO.DOC)
-- DECLARA��O DE VARI�VEL INTEIRA NA ENTIDADE PRINCIPAL

ENTITY PROJETO05 IS
PORT ( A : IN INTEGER RANGE 0 TO 7 ;
       S : OUT BIT               ) ;
END PROJETO05 ;

ARCHITECTURE PROJ05 OF PROJETO05 IS
BEGIN

WITH A SELECT
S <= '1' WHEN 0 ,
     '0' WHEN 1 ,
     '1' WHEN 2 ,
     '1' WHEN 3 ,
     '1' WHEN 4 ,
     '0' WHEN 5 ,
     '1' WHEN 6 ,
     '0' WHEN 7 ;
     
END PROJ05 ;