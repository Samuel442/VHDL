
-- IMPLEMENTA��O DE UM DEMULTIPLEXADOR 1x4 CONFORME CIRCUITO 03 DO ARQUIVO ANEXO (COMPLEMENTO.DOC)
-- DECLARA��O DE VARI�VEL INTEIRA NA ENTIDADE PRINCIPAL

ENTITY PROJETO08 IS
PORT ( E : IN BIT                  ; 
       A : IN INTEGER RANGE 0 TO 3 ;
       S0, S1, S2, S3 : OUT BIT  ) ;
END PROJETO08 ;

ARCHITECTURE PROJ08 OF PROJETO08 IS
BEGIN

S0 <= E WHEN A = 0 ELSE '1' ;
S1 <= E WHEN A = 1 ELSE '1' ;
S2 <= E WHEN A = 2 ELSE '1' ;
S3 <= E WHEN A = 3 ELSE '1' ;
     
END PROJ08 ;