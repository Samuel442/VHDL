
-- CONTADOR S�NCRONO DE D�CADA (CIRCUITO 10) DO ARQUIVO ANEXO (COMPLEMENTO.DOC)

ENTITY PROJETO16 IS
PORT ( CLOCK, CLEAR : IN BIT ;
	   QOUT         : BUFFER BIT_VECTOR (3 DOWNTO 0));
END PROJETO16 ;

ARCHITECTURE PROJ16 OF PROJETO16 IS

	COMPONENT PROJETO12
	PORT (PRN, CLRN, CLKN, J, K : IN BIT;
      Q : BUFFER BIT ) ;
	END COMPONENT; 

BEGIN

FF0: PROJETO12 PORT MAP( J => '1',                                   K => '1',                 PRN => '1', CLRN => CLEAR, CLKN => CLOCK, Q => QOUT(0) );
FF1: PROJETO12 PORT MAP( J => QOUT(0) AND (NOT QOUT(3)),             K => QOUT(0),             PRN => '1', CLRN => CLEAR, CLKN => CLOCK, Q => QOUT(1) );
FF2: PROJETO12 PORT MAP( J => QOUT(1) AND QOUT(0),                   K => QOUT(1) AND QOUT(0), PRN => '1', CLRN => CLEAR, CLKN => CLOCK, Q => QOUT(2) );
FF3: PROJETO12 PORT MAP( J => QOUT(2) AND QOUT(1) AND QOUT(0),       K => QOUT(0),             PRN => '1', CLRN => CLEAR, CLKN => CLOCK, Q => QOUT(3) );

END PROJ16;


-- COMPONENTE: FLIP FLOP JK MESTRE ESCRAVO COM PRESET E CLEAR

ENTITY PROJETO12 IS
PORT (PRN, CLRN, CLKN, J, K : IN BIT;
      Q : BUFFER BIT ) ;
END PROJETO12 ;

ARCHITECTURE PROJ12 OF PROJETO12 IS

BEGIN

PROCESS ( PRN, CLRN, CLKN )
	BEGIN
		IF     PRN = '0' THEN Q <= '1' ;
		ELSIF CLRN = '0' THEN Q <= '0' ;
		ELSIF CLKN = '0' AND CLKN 'EVENT THEN 
			IF    J = '1' AND K = '1' THEN Q <= NOT Q ;
		    ELSIF J = '1' AND K = '0' THEN Q <= '1' ;
		    ELSIF J = '0' AND K = '1' THEN Q <= '0' ;
			END IF ;
		END IF;
	END PROCESS ;
	Q <= Q ;
END PROJ12 ;
